module top;
  initial begin
    $display("HELLO, World");
    $finish;
  end
endmodule
